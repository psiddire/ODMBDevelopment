
// file: ibert_ultrascale_gth_0.v
//////////////////////////////////////////////////////////////////////////////
//   ____  ____
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 2012.3
//  \   \         Application : IBERT 7Series
//  /   /         Filename : example_ibert_ultrascale_gth_0
// /___/   /\
// \   \  /  \
//  \___\/\___\
//
//
// Module example_ibert_ultrascale_gth_0
// Generated by Xilinx IBERT_7S
//////////////////////////////////////////////////////////////////////////////

`define C_NUM_GTH_QUADS 1
`define C_GTH_REFCLKS_USED 1
module example_ibert_ultrascale_gth_0
(
  // GT top level ports
  output [(4*`C_NUM_GTH_QUADS)-1:0]     DAQ_TX_N,
  output [(4*`C_NUM_GTH_QUADS)-1:0]	    DAQ_TX_P,
  input  [(4*`C_NUM_GTH_QUADS)-1:1]    	B04_RX_N,
  input  [(4*`C_NUM_GTH_QUADS)-1:1]   	B04_RX_P,
  input                                 BCK_PRS_N,
  input                                 BCK_PRS_P,
  input                           	    GP_CLK_6_P,
  input                           	    GP_CLK_6_N,
  input  [`C_GTH_REFCLKS_USED-1:0]      REF_CLK_2_P,
  input  [`C_GTH_REFCLKS_USED-1:0]      REF_CLK_2_N,
  input  [`C_GTH_REFCLKS_USED-1:0]      REF_CLK_5_P,
  input  [`C_GTH_REFCLKS_USED-1:0]      REF_CLK_5_N,
  output                                B04_I2C_ENA,
  output                                B04_CS_B,
  output                                B04_RST_B,
  output                                KUS_DL_SEL,
  output                                FPGA_SEL,
  output                                RST_CLKS_B
);

  //
  // Ibert refclk internal signals
  //
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk1_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk1_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk1_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk11_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk11_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk11_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_refclk0_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_refclk1_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_odiv2_0_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_odiv2_1_i;
  wire                            gth_sysclk_i;
  wire   		            	  clk_gp6;

  wire  [(4*`C_NUM_GTH_QUADS)-1:0] gth_txn_o;
  wire  [(4*`C_NUM_GTH_QUADS)-1:0] gth_txp_o;
  wire  [(4*`C_NUM_GTH_QUADS)-1:0] gth_rxn_i;
  wire  [(4*`C_NUM_GTH_QUADS)-1:0] gth_rxp_i;

  // Constant driver for selector/reset pins for board to work
  assign KUS_DL_SEL = 1'b1;
  assign FPGA_SEL = 1'b0;
  assign RST_CLKS_B = 1'b1;

  // Constant driver for firefly selector/reset pins
  assign B04_I2C_ENA = 1'b0;
  assign B04_CS_B = 1'b1;
  assign B04_RST_B = 1'b1;

  // Quad 227 <-- there should be at least 1 quad
  assign gth_rxp_i[0] = BCK_PRS_P;
  assign gth_rxn_i[0] = BCK_PRS_N;
  assign gth_rxp_i[(4*`C_NUM_GTH_QUADS)-1:1] = B04_RX_P;
  assign gth_rxn_i[(4*`C_NUM_GTH_QUADS)-1:1] = B04_RX_N;

  assign DAQ_TX_P = gth_txp_o;
  assign DAQ_TX_N = gth_txn_o;

  //
  // Refclk IBUFDS instantiations
  //
    IBUFDS_GTE3 u_buf_gth_q3_clk0
      (
        .O            (gth_refclk0_i[0]),
        .ODIV2        (gth_odiv2_0_i[0]),
        .CEB          (1'b0),
        .I            (REF_CLK_2_P[0]),
        .IB           (REF_CLK_2_N[0])
      );

    IBUFDS_GTE3 u_buf_gth_q3_clk1
      (
        .O            (gth_refclk1_i[0]),
        .ODIV2        (gth_odiv2_1_i[0]),
        .CEB          (1'b0),
        .I            (REF_CLK_5_P[0]),
        .IB           (REF_CLK_5_N[0])
      );

  //
  // Refclk connection from each IBUFDS to respective quads depending on the source selected in gui
  //
  assign gth_qrefclk0_i[0] = gth_refclk0_i[0];
  assign gth_qrefclk1_i[0] = gth_refclk1_i[0];
  assign gth_qnorthrefclk0_i[0] = 1'b0;
  assign gth_qnorthrefclk1_i[0] = 1'b0;
  assign gth_qsouthrefclk0_i[0] = 1'b0;
  assign gth_qsouthrefclk1_i[0] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[0] = gth_refclk0_i[0];
  assign gth_qrefclk10_i[0] = gth_refclk1_i[0];
  assign gth_qrefclk01_i[0] = 1'b0;
  assign gth_qrefclk11_i[0] = 1'b0;
  assign gth_qnorthrefclk00_i[0] = 1'b0;
  assign gth_qnorthrefclk10_i[0] = 1'b0;
  assign gth_qnorthrefclk01_i[0] = 1'b0;
  assign gth_qnorthrefclk11_i[0] = 1'b0;
  assign gth_qsouthrefclk00_i[0] = 1'b0;
  assign gth_qsouthrefclk10_i[0] = 1'b0;
  assign gth_qsouthrefclk01_i[0] = 1'b0;
  assign gth_qsouthrefclk11_i[0] = 1'b0;


  //
  // Sysclock IBUFDS instantiation
  //
  IBUFGDS
   #(.DIFF_TERM("FALSE"))
   u_ibufgds
    (
      .I(GP_CLK_6_P),
      .IB(GP_CLK_6_N),
      .O(clk_gp6)
    );

  // Adding BUFG to the clocks
  BUFG
   u_bufg_gp6
    (
      .I(clk_gp6),
      .O(gth_sysclk_i)
    );

  //
  // IBERT core instantiation
  //
  ibert_ultrascale_gth_0 u_ibert_gth_core
    (
      .txn_o(gth_txn_o),
      .txp_o(gth_txp_o),
      .rxn_i(gth_rxn_i),
      .rxp_i(gth_rxp_i),
      .clk(gth_sysclk_i),
      .gtrefclk0_i(gth_qrefclk0_i),
      .gtrefclk1_i(gth_qrefclk1_i),
      .gtnorthrefclk0_i(gth_qnorthrefclk0_i),
      .gtnorthrefclk1_i(gth_qnorthrefclk1_i),
      .gtsouthrefclk0_i(gth_qsouthrefclk0_i),
      .gtsouthrefclk1_i(gth_qsouthrefclk1_i),
      .gtrefclk00_i(gth_qrefclk00_i),
      .gtrefclk10_i(gth_qrefclk10_i),
      .gtrefclk01_i(gth_qrefclk01_i),
      .gtrefclk11_i(gth_qrefclk11_i),
      .gtnorthrefclk00_i(gth_qnorthrefclk00_i),
      .gtnorthrefclk10_i(gth_qnorthrefclk10_i),
      .gtnorthrefclk01_i(gth_qnorthrefclk01_i),
      .gtnorthrefclk11_i(gth_qnorthrefclk11_i),
      .gtsouthrefclk00_i(gth_qsouthrefclk00_i),
      .gtsouthrefclk10_i(gth_qsouthrefclk10_i),
      .gtsouthrefclk01_i(gth_qsouthrefclk01_i),
      .gtsouthrefclk11_i(gth_qsouthrefclk11_i)
    );

endmodule
